module top_module( input in, output out );
    not ( out, in);
endmodule
